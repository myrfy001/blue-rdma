import DataTypes :: *;

typedef 0 USER_LOGIC_XDMA_TUSER_WIDTH;
typedef 512 USER_LOGIC_XDMA_DATA_WIDTH;
typedef TDiv#(USER_LOGIC_XDMA_DATA_WIDTH, 8) USER_LOGIC_XDMA_KEEP_WIDTH;

// Make sure USER_LOGIC_DESCRIPTOR_BIT_WIDTH * USER_LOGIC_RING_BUF_DEEP = 4kB
typedef 32   USER_LOGIC_DESCRIPTOR_BYTE_WIDTH;
typedef TMul#(USER_LOGIC_DESCRIPTOR_BYTE_WIDTH, BYTE_WIDTH)  USER_LOGIC_DESCRIPTOR_BIT_WIDTH; // 256 bit
typedef 128  USER_LOGIC_RING_BUF_DEEP; 
typedef TLog#(USER_LOGIC_RING_BUF_DEEP)  USER_LOGIC_RING_BUF_DEEP_WIDTH ; 



typedef 2 RINGBUF_H2C_TOTAL_COUNT;
typedef 2 RINGBUF_C2H_TOTAL_COUNT;

typedef 3 RINGBUF_NUMBER_WIDTH;


typedef 4 CSR_DATA_BYTE_NUM;
typedef TLog#(CSR_DATA_BYTE_NUM) CSR_ADDR_INTERVAL_WIDTH;  // 2 bit
typedef 1048576 PCIE_CONFIG_BAR_SPACE_BYTE_SIZE;  // 1024 * 1024
typedef TLog#(PCIE_CONFIG_BAR_SPACE_BYTE_SIZE) PCIE_CONFIG_BAR_SPACE_BYTE_WIDTH;

// CSR are grouped into 4kB groups, each CSR is 4 bytes width, so each group has 1024 entry.
typedef 1024 CSR_GROUP_ENTRY_CNT;
typedef TLog#(CSR_GROUP_ENTRY_CNT) CSR_GROUP_WIDTH;

// how many CSR groups can the config BAR space hold.
typedef TSub#(PCIE_CONFIG_BAR_SPACE_BYTE_WIDTH, TAdd#(CSR_ADDR_INTERVAL_WIDTH, CSR_GROUP_WIDTH)) CSR_GROUP_CNT_WIDTH;





typedef 16 CMD_QUEUE_DESCRIPTOR_MAX_SEGMENT_CNT;

typedef 2024042901 HARDWARE_VERSION;