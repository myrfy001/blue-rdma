typedef 0 USER_LOGIC_XDMA_TUSER_WIDTH;
typedef 256 USER_LOGIC_XDMA_DATA_WIDTH;
typedef TDiv#(USER_LOGIC_XDMA_DATA_WIDTH, 8) USER_LOGIC_XDMA_KEEP_WIDTH;