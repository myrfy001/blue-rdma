import RdmaUtils :: *;

import QPContext :: *;

(* doc = "testcase" *)
module mkTestQueryContxt(Empty);
    
endmodule