import ClientServer :: *;
import GetPut :: *;

import DataTypes :: *;
import UserLogicSettings :: *;

interface CommandQueueController;
    
endinterface