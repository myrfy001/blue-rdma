import RQ :: *;

(* doc = "testcase" *)
module mkTestRqQueryContxt(Empty);
    
endmodule