typedef 0 USER_LOGIC_XDMA_TUSER_WIDTH;
typedef 256 USER_LOGIC_XDMA_DATA_WIDTH;
typedef TDiv#(USER_LOGIC_XDMA_DATA_WIDTH, 8) USER_LOGIC_XDMA_KEEP_WIDTH;

// Make sure USER_LOGIC_DESCRIPTOR_BIT_WIDTH * USER_LOGIC_RING_BUF_LEN = 4kB
typedef 32   USER_LOGIC_DESCRIPTOR_BYTE_WIDTH;
typedef TMul#(USER_LOGIC_DESCRIPTOR_BYTE_WIDTH, BYTE_WIDTH)  USER_LOGIC_DESCRIPTOR_BIT_WIDTH; // 256 bit
typedef 128  USER_LOGIC_RING_BUF_LEN; 
typedef TLog#(USER_LOGIC_RING_BUF_LEN)  USER_LOGIC_RING_BUF_LEN_WIDTH ; 


typedef 2 RINGBUF_H2C_TOTAL_COUNT;
typedef 2 RINGBUF_C2H_TOTAL_COUNT;
typedef TAdd#(RINGBUF_H2C_TOTAL_COUNT, RINGBUF_C2H_TOTAL_COUNT) RINGBUF_TOTAL_COUNT;
typedef TLog#(RINGBUF_TOTAL_COUNT) RINGBUF_INDEX_WIDTH;
typedef Bit#(RINGBUF_INDEX_WIDTH) RingbufIndex;
